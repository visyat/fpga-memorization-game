module display();

endmodule